module ConditionCheck();






endmodule
