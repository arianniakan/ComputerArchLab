module ControlUnit(input S, input mode [1:0], input Op-code [3:0], output Execute_Command [3:0],
                   output mem_read, output mem_write,output WB_enable,output B,output Status_Reg_Update);





















endmodule