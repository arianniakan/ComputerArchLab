module arm(input clk, rst);
endmodule