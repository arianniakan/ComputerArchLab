module ARM_DP_tb;
reg clk;
reg rst_n;

 
ARM_DP uut(
    .rst (rst_n),
    .clk (clk)
);

localparam CLK_PERIOD = 10;
always #(CLK_PERIOD/2) clk=~clk;

initial begin
    #1 rst_n<=1'bx;clk<=1'bx;
    #(CLK_PERIOD*3) rst_n<=1;
    #(CLK_PERIOD*3) rst_n<=0;clk<=0;
    repeat(5) @(posedge clk);
    @(posedge clk);
    repeat(2) @(posedge clk);
    #1000 $stop;
end

endmodule
