module RegisterFile( input clk, rst, input [3:0] src1, src2, Dest_eb, 
                    input [31:0] Result_WB, 
                    input writeBackEn, 
                    output [31:0] reg1, reg2);
reg [31:0] REGISTERS [0:16];



endmodule