module ConditionCheck()