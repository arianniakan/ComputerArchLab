module ControlUnit (input S, input [1:0]  mode, input [3:0] Op_code, output [3:0] Execute_Command,
                   output mem_read, output mem_write,output WB_enable, output B, output Status_Reg);


endmodule